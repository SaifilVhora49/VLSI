module mux8x1_tb;
	reg[2:0] s;
	reg[7:0] in;
	wire out;
	mux8x1 uut(in,s,out);
	initial begin
	s[0]=0; s[1]=0; s[2]=0; in[0]=0; in[1]=0; in[2]=0;in[3]=0;in[4]=0;in[5]=0;in[6]=0;in[7]=0;
	#10 in[0]=1;
	#10 s[0]=1;
	#10 in[1]=1;
	#10 s[1]=1; s[0]=0;
	#10 in[2]=1;
	#10 s[1]=1; s[0]=1;
	#10 in[3]=1;
	#10 s[1]=0; s[0]=0; s[2]=1;
	#10 in[4]=1;
	#10 s[1]=1; s[0]=0; s[2]=1;
	#10 in[5]=1;
	#10 s[1]=0; s[0]=1; s[2]=1;
	#10 in[6]=1;
	#10 s[1]=1; s[0]=1; s[2]=1;
	end
endmodule
	
